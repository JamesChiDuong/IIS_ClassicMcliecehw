
module Data_Transmitter(
    input clk,                                          
    output o_uart_tx
    );
localparam  DBITS = 8,                              // 8 bit data
            BR_LIMIT = 53,                          // counter limit value
            BR_BITS = 6,                            // number of counter bits
            SB_TICK = 16,
            WELCOME_STR_LEN = 21;                   // String lengh of the Welcom string   
reg [DBITS-1:0] WELCOME_STR[0:WELCOME_STR_LEN-1];   // Init array Data
reg [4:0] tx_index = 0;                             // the index of the String
wire tx_done;                                       // Check when the transfer data done
reg tx_Send;                                        // Start to send the Data
reg [DBITS-1:0] tx_data = 0;                        // Buffer Data
reg reset;                                          // Reset signal
wire tick;                                          // Tick signal which is generated by baudate




/***********Initilation the String "Hello world******************/
reg [27:0] counter;
initial begin
    WELCOME_STR[1]   = "H";
    WELCOME_STR[2]   = "e";
    WELCOME_STR[3]   = "l";
    WELCOME_STR[4]   = "l";
    WELCOME_STR[5]   = "o";
    WELCOME_STR[6]   = " ";
    WELCOME_STR[7]   = "W";
    WELCOME_STR[8]   = "o";
    WELCOME_STR[9]   = "r";
    WELCOME_STR[10]  = "l";
    WELCOME_STR[11]  = "d";
    WELCOME_STR[12]  = " ";
    WELCOME_STR[13]  = "\r";
    WELCOME_STR[14]  = "\n";
end

// assign tx_fifo_not_empty = ~tx_empty;
initial counter = 28'hffffff0;
initial tx_index = 5'd0;
initial tx_Send = 1'b0;
initial	reset = 1'b1;
always @(posedge clk)
    reset <= 1'b0;

always @(posedge clk) begin
    counter <= counter + 1'b1;                      // Counter will counter when having the clk                      
end

always @(posedge clk) begin
    if((tx_Send)&&(tx_done))                        // if the transfer finish the data and done for the transfer signal, we keep continue to transfer the next data
        tx_index <= tx_index + 1'b1;                
end

always @(posedge clk) begin                         // Assign the 1 byte data to the tx_data
    tx_data <= WELCOME_STR[tx_index];
end

always @(posedge clk) begin
    if(counter == 28'hfffffff)                      // If counter == the initial counter, it will be send the data
        tx_Send <= 1'b1;
    else if((tx_Send) && (tx_done) && (tx_index) == 5'hff)
        tx_Send <= 1'b0;                            // If transfer done,signal tx_send =1 and the full of the string welcome is reached, it will stop
end
baud_rate_generator 
    #(
        .N(BR_BITS), 
        .M(BR_LIMIT)
     ) 
    BAUD_RATE_GEN   
    (
        .clk(clk), 
        .reset(reset),
        .tick(tick)
     );

Transmitter
    #(
        .DBITS(DBITS),
        .SB_TICK(SB_TICK)
     )
     UART_TX_UNIT
     (
        .clk(clk),
        .reset(reset),
        .tx_start(tx_Send),
        .sample_tick(tick),
        .data_in(tx_data),
        .tx_done(tx_done),
        .tx(o_uart_tx)
     );
endmodule